module and (A, B, out);
input A, B;

output out;

assign out = A & B;
    
endmodule